module counter(
	input wire clk,
	input wire rst_n,
	output wire [9:0] cnt
);

reg [9:0] cnt_r;

always @(posedge clk or negedge rst_n)
	if (rst_n == 1'b0)
		cnt_r <= 10'd0;
	else
		cnt_r = cnt_r + 1'b1;
		
assign cnt = cnt_r;

endmodule